library IEEE;
use IEEE.std_logic_1164.all;
--- entity declaration
entity NOT_1 is
	port(I0 : in std_logic;
		  O0 : out std_logic);
end entity;

architecture functionality of NOT_1 is

begin
	O0 <= NOT I0;
end functionality;
