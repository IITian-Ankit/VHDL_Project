library IEEE;
use 